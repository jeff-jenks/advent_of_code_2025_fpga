`define ASCII_EOT 8'h04 // End of Transmission
`define ASCII_LF 8'h0A // Line Feed
`define ASCII_NUM 8'h23 // # Number Sign
`define ASCII_CLOSE_PAR 8'h29 // ) Close parenthesis
`define ASCII_PERIOD 8'h2E // . Period
`define ASCII_0 8'h30 // 0 Zero
`define ASCII_1 8'h31 // 1 One
`define ASCII_2 8'h32 // 2 Two
`define ASCII_3 8'h33 // 3 Three
`define ASCII_4 8'h34 // 4 Four
`define ASCII_5 8'h35 // 5 Five
`define ASCII_6 8'h36 // 6 Six
`define ASCII_7 8'h37 // 7 Seven
`define ASCII_8 8'h38 // 8 Eight
`define ASCII_9 8'h39 // 9 Nine
`define ASCII_F 8'h46 // F Capital F
`define ASCII_P 8'h50 // P Capital P
`define ASCII_S 8'h53 // S Capital S
`define ASCII_CARET 8'h5E // ^ Caret
`define ASCII_OPEN_BRACE 8'h7B // { Opening brace
`define ASCII_CLOSE_BRACE 8'h7D // } Closing brace
